
`define BLIT_NOP  5'd0
`define BLIT_RECT 5'd1
`define BLIT_COPY 5'd2
`define BLIT_TEXT 5'd3
